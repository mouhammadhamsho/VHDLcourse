library verilog;
use verilog.vl_types.all;
entity ProgramCounterTopLevel_vlg_vec_tst is
end ProgramCounterTopLevel_vlg_vec_tst;
