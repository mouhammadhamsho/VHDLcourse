library ieee;
use ieee.std_logic_1164.all;

entity SR_Latch_EN is

generic(
N : Integer := 8);


port(
S , R,EN : in std_logic;
Q, QN : out std_logic

);
end  SR_Latch_EN;

architecture behavioral of SR_Latch_EN is 


signal Q_temp , QN_temp : std_logic;

begin

Q_temp<=(R AND EN) NOR QN_temp;
QN_temp<= (S AND EN) NOR Q_temp;


Q<=Q_temp;
QN<=QN_temp;

end;
 