library verilog;
use verilog.vl_types.all;
entity ModulePCRAM_vlg_vec_tst is
end ModulePCRAM_vlg_vec_tst;
