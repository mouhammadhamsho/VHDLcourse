library verilog;
use verilog.vl_types.all;
entity ProgramCounterTopLevel_vlg_check_tst is
    port(
        PC_COUNT_OUT    : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end ProgramCounterTopLevel_vlg_check_tst;
